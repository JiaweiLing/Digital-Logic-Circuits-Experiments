`timescale 10 ns/ 1 ps
module test_decode416(); 
reg [3:0] x;
reg en; 
wire [15:0]y;
decode416 i1( .x(x),.en(en),.y(y));

initial begin
en =1’b1; x =4'b0000; #10;
		  x =4'b0001; #10;
		  x =4'b0010; #10;
		  x =4'b0011; #10;
		  x =4'b0100; #10;
		  x =4'b0101; #10;
		  x =4'b0110; #10;
		  x =4'b0111; #10;
		  x =4'b1000; #10;
		  x =4'b1001; #10;
		  x =4'b1010; #10;
		  x =4'b1011; #10;
		  x =4'b1100; #10;
		  x =4'b1101; #10;
		  x =4'b1110; #10;
		  x =4'b1111; #10;
en =1’b0; x =4'b0000; #10;
		  x =4'b0001; #10;
		  x =4'b0010; #10;
		  x =4'b0011; #10;
		  x =4'b0100; #10;
		  x =4'b0101; #10;
		  x =4'b0110; #10;
		  x =4'b0111; #10;
		  x =4'b1000; #10;
		  x =4'b1001; #10;
		  x =4'b1010; #10;
		  x =4'b1011; #10;
		  x =4'b1100; #10;
		  x =4'b1101; #10;
		  x =4'b1110; #10;
		  x =4'b1111; #10;
	end
endmodule